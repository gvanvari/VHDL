library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.std_logic_unsigned.all;

entity input_ROM is
PORT (
    i: IN STD_LOGIC_VECTOR(4 downto 0);
    inp_sel: IN STD_LOGIC_VECTOR(1 downto 0);
    o_r: OUT STD_LOGIC_VECTOR(31 downto 0);
    o_i: OUT STD_LOGIC_VECTOR(31 downto 0));
end input_ROM;

architecture Behavioral of input_ROM is
TYPE marray is array(0 to 31) of std_logic_vector(31 downto 0);
CONSTANT real1 : marray:=(X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000");
CONSTANT imag1 : marray:=(X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000",X"3f800000");
CONSTANT real2 : marray:=(X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000");
CONSTANT imag2 : marray:=(X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000",X"40000000");
CONSTANT real3 : marray:=(X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000");
CONSTANT imag3 : marray:=(X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000",X"40400000");
CONSTANT real4 : marray:=(X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000");
CONSTANT imag4 : marray:=(X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000",X"40800000");

begin
with inp_sel select
o_r <= real1(conv_integer(i)) when "00",
real2(conv_integer(i)) when "01",
real3(conv_integer(i)) when "10",
real4(conv_integer(i)) when others;

with inp_sel select
o_i <= imag1(conv_integer(i)) when "00",
imag2(conv_integer(i)) when "01",
imag3(conv_integer(i)) when "10",
imag4(conv_integer(i)) when others;
end Behavioral;
